  
class DataCtrl;
  // Declare four logic 8-bit wide class attributes. Name attributes data1, data2, data3, data4
  logic [7:0] data1, data2, data3, data4;
  
endclass